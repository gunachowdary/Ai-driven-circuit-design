* Simple RC Circuit
V1 1 0 DC 5
R1 1 2 1k
C1 2 0 1u
.tran 0.1ms 10ms UIC
.ic v(2) = 0
.plot tran v(2)
.end
